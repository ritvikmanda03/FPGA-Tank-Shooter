module finalbullet_rom (
	input logic clock,
	input logic [5:0] address,
	output logic [3:0] q
);

logic [3:0] memory [0:48] /* synthesis ram_init_file = "./finalbullet/finalbullet.mif" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
