module floor2_rom (
	input logic clock,
	input logic [14:0] address,
	output logic [3:0] q
);

logic [3:0] memory [0:20479] /* synthesis ram_init_file = "./floor2/floor2.mif" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
